/******************************************************************************

File name:    initiator_bram.v
Rev:          5.4
Description:  This is the Initiator BRAM (IRAM) module of the
              User Design. It stores preloaded field information
              with different data patterns. This data is used to 
              populate the DATA field of outgoing Initiator Request 
              packets from the IREQ Generator module. The IRAM is 
              also used by the IRESP Handler to verify the DATA 
              field of incoming Initiator Response packets against 
              the expected contents.

#-- Copyright (c) 1995-2008 by Xilinx, Inc. All rights reserved.
#-- This text/file contains proprietary, confidential
#-- information of Xilinx, Inc., is distributed under license
#-- from Xilinx, Inc., and may be used, copied and/or
#-- disclosed only pursuant to the terms of a valid license
#-- agreement with Xilinx, Inc. Xilinx hereby grants you a
#-- license to use this text/file solely for design, simulation,
#-- implementation and creation of design files limited
#-- to Xilinx devices or technologies. Use with non-Xilinx
#-- devices or technologies is expressly prohibited and
#-- immediately terminates your license unless covered by
#-- a separate agreement.
#--
#-- Xilinx is providing this design, code, or information
#-- "as-is" solely for use in developing programs and
#-- solutions for Xilinx devices, with no obligation on the
#-- part of Xilinx to provide support. By providing this design,
#-- code, or information as one possible implementation of
#-- this feature, application or standard, Xilinx is making no
#-- representation that this implementation is free from any
#-- claims of infringement. You are responsible for
#-- obtaining any rights you may require for your implementation.
#-- Xilinx expressly disclaims any warranty whatsoever with
#-- respect to the adequacy of the implementation, including
#-- but not limited to any warranties or representations that this
#-- implementation is free from claims of infringement, implied
#-- warranties of merchantability or fitness for a particular
#-- purpose.
#--
#-- Xilinx products are not intended for use in life support
#-- appliances, devices, or systems. Use in such applications is
#-- expressly prohibited.
#--
#-- Any modifications that are made to the Source Code are
#-- done at the user's sole risk and will be unsupported.
#--
#-- This copyright and support notice must be retained as part
#-- of this text at all times. (c) Copyright 1995-2008 Xilinx, Inc.
#-- All rights reserved.
*******************************************************************************/
`timescale 1 ps / 1 ps

module initiator_bram #(
  parameter TCQ = 100
)(

  // System
  input           lnk_clk,      // Link clock
  input           lnk_reset_n,  // Active low reset

  // IREQ Generator
  input   [0:9]   g_iram_addra, // Address from IREQ Generator into IRAM
  output  [0:63]  iram_doa,     // Read data from IRAM to IREQ Generator

  // IRESP Handler
  input   [0:9]   h_iram_addrb, // Address from IRESP Handler into IRAM
  output  [0:63]  iram_dob      // Read data from IRAM to IRESP Handler
  );

  // Construct Initiator BRAM from two 1kx36 RAMB36 primitives cascaded in 
  // width resulting in a 1kx64 memory. The IRAM wil be put into WRITE_FIRST
  // mode to allow for a write path to be added from the Bypass Port. 
  //
  // The IRAM will be initialized with the following data patterns:
  //
  // Address Range  |   Data Type 
  // -------------------------------------------------------
  // 0x000 - 0x01F  |   All 0�s
  // 0x020 - 0x03F  |   All 1�s
  // 0x040 - 0x05F  |   Alternating 0�s and 1�s
  // 0x060 - 0x07F  |   Alternating 1�s and 0�s
  // 0x080 - 0x09F  |   Alternating bytes of 0�s and 1�s
  // 0x0A0 - 0x0BF  |   Alternating bytes of 1�s and 0�s
  // 0x0C0 - 0x0DF  |   Alternating dwords of 0�s and 1�s
  // 0x0E0 - 0x0FF  |   Alternating dwords of 1�s and 0�s
  // 0x100 - 0x11F  |   Incrementing bytes
  // 0x120 - 0x13F  |   Incrementing dwords
  // 0x140 - 0x15F  |   Decrementing bytes
  // 0x160 - 0x17F  |   Decrementing dwords
  // 0x180 - 0x19F  |   Random data #1
  // 0x1A0 - 0x1BF  |   Random data #2
  // 0x1C0 - 0x7FF  |   More incrementing dwords
  
  RAMB36 #(
    .READ_WIDTH_A(36),
    .READ_WIDTH_B(36),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(36),
    .WRITE_WIDTH_B(36),
    // The following INIT_xx declarations specify the initial contents of the RAM.
    // These INITs specify the lower 32 bits of the pattern. The INITs of the other
    // BRAM initialize the upper 32 bits of the pattern.
    // All 0's
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    // All 1's
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    // Alternating 0's and 1's
    .INIT_08(256'h5555555555555555555555555555555555555555555555555555555555555555),
    .INIT_09(256'h5555555555555555555555555555555555555555555555555555555555555555),
    .INIT_0A(256'h5555555555555555555555555555555555555555555555555555555555555555),
    .INIT_0B(256'h5555555555555555555555555555555555555555555555555555555555555555),
    // Alternating 1's and 0's
    .INIT_0C(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_0D(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_0E(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_0F(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    // Alternating bytes of 0's and 1's
    .INIT_10(256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF),
    .INIT_11(256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF),
    .INIT_12(256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF),
    .INIT_13(256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF),
    // Alternating bytes of 1's and 0's
    .INIT_14(256'hFF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00),
    .INIT_15(256'hFF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00),
    .INIT_16(256'hFF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00),
    .INIT_17(256'hFF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00),
    // Alternating dwords of 0's and 1's
    .INIT_18(256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF),
    .INIT_19(256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF),
    .INIT_1A(256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF),
    .INIT_1B(256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF),
    // Alternating dwords of 1's and 0's
    .INIT_1C(256'hFFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000),
    .INIT_1D(256'hFFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000),
    .INIT_1E(256'hFFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000),
    .INIT_1F(256'hFFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000),
    // Incrementing bytes
    .INIT_20(256'h0001020308090A0B1011121318191A1B2021222328292A2B3031323338393A3B),
    .INIT_21(256'h4041424348494A4B5051525358595A5B6061626368696A6B7071727378797A7B),
    .INIT_22(256'h8081828388898A8B9091929398999A9BA0A1A2A3A8A9AAABB0B1B2B3B8B9BABB),
    .INIT_23(256'hC0C1C2C3C8C9CACBD0D1D2D3D8D9DADBE0E1E2E3E8E9EAEBF0F1F2F3F8F9FAFB),
    // Incrementing dwords
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    // Decrementing bytes
    .INIT_28(256'hFFFEFDFCF7F6F5F4EFEEEDECE7E6E5E4DFDEDDDCD7D6D5D4CFCECDCCC7C6C5C4),
    .INIT_29(256'hBFBEBDBCB7B6B5B4AFAEADACA7A6A5A49F9E9D9C979695948F8E8D8C87868584),
    .INIT_2A(256'h7F7E7D7C777675746F6E6D6C676665645F5E5D5C575655544F4E4D4C47464544),
    .INIT_2B(256'h3F3E3D3C373635342F2E2D2C272625241F1E1D1C171615140F0E0D0C07060504),
    // Decrementing dwords
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    // Random Data #1
    .INIT_30(256'h40888BA10E82FB03102131AA6A65B7048B2927D64F4B4A3102131AA6A645ACFD),
    .INIT_31(256'h7AD9B0660014D920876D1A3C3864C04A63FD41FF1BB79B4A310F7B7BB8F5D24A),
    .INIT_32(256'h2B6A923ED08B8920E5CFEC97EB7015209C9EEE8D14C70480F69A24C1916C4880),
    .INIT_33(256'hF9F973DFA353BC80AC3EBE1D53BA14801A355FDFED38C3004482EF8D40A54300),
    // Random Data #2
    .INIT_34(256'hFC28767E796E3800C93D200EAE38D0007CE423368056D00094935192586A1321),
    .INIT_35(256'hE44049B62503D656E60909F7F2073031640611E4D37B8F3B2DCA845E70AF3171),
    .INIT_36(256'hC0E5C09F37CE6792E479B612E12A10A548D99E92943DFE47F3989BF6972EAA49),
    .INIT_37(256'h72497F5F50DCA3A8C03F35E38192F028680F84CDE62FB1B0576AB47AED8622B0),
    // More incrementing dwords
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000)

    ) iram_upper (
    .DOA(iram_doa[0:31]),
    .DOB(iram_dob[0:31]),
    .DOPA( ),
    .DOPB( ),
    .ADDRA({1'b0, g_iram_addra, 5'b0}),
    .ADDRB({1'b0, h_iram_addrb, 5'b0}),
    .CLKA(lnk_clk),
    .CLKB(lnk_clk),
    .DIA(32'b0),
    .DIB(32'b0),
    .DIPA(4'b0),
    .DIPB(4'b0),
    .ENA(1'b1),
    .ENB(1'b1),
    .REGCEA(1'b0),
    .REGCEB(1'b0),
    .SSRA(~lnk_reset_n),
    .SSRB(~lnk_reset_n),
    .WEA(4'b0),
    .WEB(4'b0),
    .CASCADEOUTLATA(),
    .CASCADEOUTLATB(),
    .CASCADEOUTREGA(),
    .CASCADEOUTREGB(),
    .CASCADEINLATA(),
    .CASCADEINLATB(),
    .CASCADEINREGA(),
    .CASCADEINREGB()
    );


  RAMB36 #(
    .READ_WIDTH_A(36),
    .READ_WIDTH_B(36),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(36),
    .WRITE_WIDTH_B(36),
    // The following INIT_xx declarations specify the initial contents of the RAM.
    // These INITs specify the lower 32 bits of the pattern. The INITs of the other
    // BRAM initialize the upper 32 bits of the pattern.
    // All 0's
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    // All 1's
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    // Alternating 0's and 1's
    .INIT_08(256'h5555555555555555555555555555555555555555555555555555555555555555),
    .INIT_09(256'h5555555555555555555555555555555555555555555555555555555555555555),
    .INIT_0A(256'h5555555555555555555555555555555555555555555555555555555555555555),
    .INIT_0B(256'h5555555555555555555555555555555555555555555555555555555555555555),
    // Alternating 1's and 0's
    .INIT_0C(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_0D(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_0E(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_0F(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    // Alternating bytes of 0's and 1's
    .INIT_10(256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF),
    .INIT_11(256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF),
    .INIT_12(256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF),
    .INIT_13(256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF),
    // Alternating bytes of 1's and 0's
    .INIT_14(256'hFF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00),
    .INIT_15(256'hFF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00),
    .INIT_16(256'hFF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00),
    .INIT_17(256'hFF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00),
    // Alternating dwords of 0's and 1's
    .INIT_18(256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF),
    .INIT_19(256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF),
    .INIT_1A(256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF),
    .INIT_1B(256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF),
    // Alternating dwords of 1's and 0's
    .INIT_1C(256'hFFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000),
    .INIT_1D(256'hFFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000),
    .INIT_1E(256'hFFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000),
    .INIT_1F(256'hFFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000),
    // Incrementing bytes
    .INIT_20(256'h040506070C0D0E0F141516171C1D1E1F242526272C2D2E2F343536373C3D3E3F),
    .INIT_21(256'h444546474C4D4E4F545556575C5D5E5F646566676C6D6E6F747576777C7D7E7F),
    .INIT_22(256'h848586878C8D8E8F949596979C9D9E9FA4A5A6A7ACADAEAFB4B5B6B7BCBDBEBF),
    .INIT_23(256'hC4C5C6C7CCCDCECFD4D5D6D7DCDDDEDFE4E5E6E7ECEDEEEFF4F5F6F7FCFDFEFF),
    // Incrementing dwords
    .INIT_24(256'h0000000000000001000000020000000300000004000000050000000600000007),
    .INIT_25(256'h00000008000000090000000A0000000B0000000C0000000D0000000E0000000F),
    .INIT_26(256'h0000001000000011000000120000001300000014000000150000001600000017),
    .INIT_27(256'h00000018000000190000001A0000001B0000001C0000001D0000001E0000001F),
    // Decrementing bytes
    .INIT_28(256'hFBFAF9F8F3F2F1E0EBEAE9E8E3E2E1E0DBDAD9D8D3D2D1D0CBCAC9C8C3C2C1C0),
    .INIT_29(256'hBBBAB9B8B3B2B1B0ABAAA9A8A3A2A1A09B9A9998939291908B8A898883828180),
    .INIT_2A(256'h7B7A7978737271706B6A6968636261605B5A5958535251504B4A494843424140),
    .INIT_2B(256'h3B3A3938333231302B2A2928232221201B1A1918131211100B0A090803020100),
    // Decrementing dwords
    .INIT_2C(256'h0000001F0000001E0000001D0000001C0000001B0000001A0000001900000018),
    .INIT_2D(256'h0000001700000016000000150000001400000013000000120000001100000010),
    .INIT_2E(256'h0000000F0000000E0000000D0000000C0000000B0000000A0000000900000008),
    .INIT_2F(256'h000000070000000600000005000000040000000B000000020000000100000000),
    // Random Data #1
    .INIT_30(256'hD2E2351827344759DFABFCDFE890AA106B7BE8C8AF9AD7E4DE7F8269906451E1),
    .INIT_31(256'h549687A4CC338D8A7D5EB4F1C3FD41FF1BB79BB6A5C156A2835D7B88D7FD5E4F),
    .INIT_32(256'hD876D1A3C3B33EEF4A42767E7ADC77D7E7F7B7BB8F5D2CC34A5D5C5DD6638710),
    .INIT_33(256'h009A54ABCDD54DD23003A102197A3EFFDFEAAB4A3102131AA6A645ACFDBBABED),
    // Random Data #2
    .INIT_34(256'hFB1CB35500555B7048B2927D64F4FAF0A95C40CFCC1B7200808373D85CB99450),
    .INIT_35(256'h81A3D3CC7DAF7B89131B3E51F16A751F55B7ED2004E501F29C2D16A6AD8F0CD4),
    .INIT_36(256'h074D9CA102C30A303864C04A6078014F8FC562376DCCDFF02240818E323B0243),
    .INIT_37(256'hC31337083756131096AF3ECAA10E013049E9A8A6121D63B03E38DEE9CDCC54D0),
    // More incrementing dwords
    .INIT_38(256'h0000000000000001000000020000000300000004000000050000000600000007),
    .INIT_39(256'h00000008000000090000000A0000000B0000000C0000000D0000000E0000000F),
    .INIT_3A(256'h0000001000000011000000120000001300000014000000150000001600000017),
    .INIT_3B(256'h00000018000000190000001A0000001B0000001C0000001D0000001E0000001F),
    .INIT_3C(256'h0000002000000021000000220000002300000024000000250000002600000027),
    .INIT_3D(256'h00000028000000290000002A0000002B0000002C0000002D0000002E0000002F),
    .INIT_3E(256'h0000003000000031000000320000003300000034000000350000003600000037),
    .INIT_3F(256'h00000038000000390000003A0000003B0000003C0000003D0000003E0000003F),
    .INIT_40(256'h0000004000000041000000420000004300000044000000450000004600000047),
    .INIT_41(256'h00000048000000490000004A0000004B0000004C0000004D0000004E0000004F),
    .INIT_42(256'h0000005000000051000000520000005300000054000000550000005600000057),
    .INIT_43(256'h00000058000000590000005A0000005B0000005C0000005D0000005E0000005F),
    .INIT_44(256'h0000006000000061000000620000006300000064000000650000006600000067),
    .INIT_45(256'h00000068000000690000006A0000006B0000006C0000006D0000006E0000006F),
    .INIT_46(256'h0000007000000071000000720000007300000074000000750000007600000077),
    .INIT_47(256'h00000078000000790000007A0000007B0000007C0000007D0000007E0000007F),
    .INIT_48(256'h0000008000000081000000820000008300000084000000850000008600000087),
    .INIT_49(256'h00000088000000890000008A0000008B0000008C0000008D0000008E0000008F),
    .INIT_4A(256'h0000009000000091000000920000009300000094000000950000009600000097),
    .INIT_4B(256'h00000098000000990000009A0000009B0000009C0000009D0000009E0000009F),
    .INIT_4C(256'h000000A0000000A1000000A2000000A3000000A4000000A5000000A6000000A7),
    .INIT_4D(256'h000000A8000000A9000000AA000000AB000000AC000000AD000000AE000000AF),
    .INIT_4E(256'h000000B0000000B1000000B2000000B3000000B4000000B5000000B6000000B7),
    .INIT_4F(256'h000000B8000000B9000000BA000000BB000000BC000000BD000000BE000000BF),
    .INIT_50(256'h000000C0000000C1000000C2000000C3000000C4000000C5000000C6000000C7),
    .INIT_51(256'h000000C8000000C9000000CA000000CB000000CC000000CD000000CE000000CF),
    .INIT_52(256'h000000D0000000D1000000D2000000D3000000D4000000D5000000D6000000D7),
    .INIT_53(256'h000000D8000000D9000000DA000000DB000000DC000000DD000000DE000000DF),
    .INIT_54(256'h000000E0000000E1000000E2000000E3000000E4000000E5000000E6000000E7),
    .INIT_55(256'h000000E8000000E9000000EA000000EB000000EC000000ED000000EE000000EF),
    .INIT_56(256'h000000F0000000F1000000F2000000F3000000F4000000F5000000F6000000F7),
    .INIT_57(256'h000000F8000000F9000000FA000000FB000000FC000000FD000000FE000000FF),
    .INIT_58(256'h0000100000000101000001020000010300000104000001050000010600000107),
    .INIT_59(256'h00001008000001090000010A0000010B0000010C0000010D0000010E0000010F),
    .INIT_5A(256'h0000101000000111000001120000011300000114000001150000011600000117),
    .INIT_5B(256'h00001018000001190000011A0000011B0000011C0000011D0000011E0000011F),
    .INIT_5C(256'h0000102000000121000001220000012300000124000001250000012600000127),
    .INIT_5D(256'h00001028000001290000012A0000012B0000012C0000012D0000012E0000012F),
    .INIT_5E(256'h0000103000000131000001320000013300000134000001350000013600000137),
    .INIT_5F(256'h00001038000001390000013A0000013B0000013C0000013D0000013E0000013F),
    .INIT_60(256'h0000104000000141000001420000014300000144000001450000014600000147),
    .INIT_61(256'h00001048000001490000014A0000014B0000014C0000014D0000014E0000014F),
    .INIT_62(256'h0000105000000151000001520000015300000154000001550000015600000157),
    .INIT_63(256'h00001058000001590000015A0000015B0000015C0000015D0000015E0000015F),
    .INIT_64(256'h0000106000000161000001620000016300000164000001650000016600000167),
    .INIT_65(256'h00001068000001690000016A0000016B0000016C0000016D0000016E0000016F),
    .INIT_66(256'h0000107000000171000001720000017300000174000001750000017600000177),
    .INIT_67(256'h00001078000001790000017A0000017B0000017C0000017D0000017E0000017F),
    .INIT_68(256'h0000108000000181000001820000018300000184000001850000018600000187),
    .INIT_69(256'h00001088000001890000018A0000018B0000018C0000018D0000018E0000018F),
    .INIT_6A(256'h0000109000000191000001920000019300000194000001950000019600000197),
    .INIT_6B(256'h00001098000001990000019A0000019B0000019C0000019D0000019E0000019F),
    .INIT_6C(256'h000010A0000001A1000001A2000001A3000001A4000001A5000001A6000001A7),
    .INIT_6D(256'h000010A8000001A9000001AA000001AB000001AC000001AD000001AE000001AF),
    .INIT_6E(256'h000010B0000001B1000001B2000001B3000001B4000001B5000001B6000001B7),
    .INIT_6F(256'h000010B8000001B9000001BA000001BB000001BC000001BD000001BE000001BF),
    .INIT_70(256'h000010C0000001C1000001C2000001C3000001C4000001C5000001C6000001C7),
    .INIT_71(256'h000010C8000001C9000001CA000001CB000001CC000001CD000001CE000001CF),
    .INIT_72(256'h000010D0000001D1000001D2000001D3000001D4000001D5000001D6000001D7),
    .INIT_73(256'h000010D8000001D9000001DA000001DB000001DC000001DD000001DE000001DF),
    .INIT_74(256'h000010E0000001E1000001E2000001E3000001E4000001E5000001E6000001E7),
    .INIT_75(256'h000010E8000001E9000001EA000001EB000001EC000001ED000001EE000001EF),
    .INIT_76(256'h000010F0000001F1000001F2000001F3000001F4000001F5000001F6000001F7),
    .INIT_77(256'h000010F8000001F9000001FA000001FB000001FC000001FD000001FE000001FF),
    .INIT_78(256'h0000200000000201000002020000020300000204000002050000020600000207),
    .INIT_79(256'h00002008000002090000020A0000020B0000020C0000020D0000020E0000020F),
    .INIT_7A(256'h0000201000000211000002120000021300000214000002150000021600000217),
    .INIT_7B(256'h00002018000002190000021A0000021B0000021C0000021D0000021E0000021F),
    .INIT_7C(256'h0000202000000221000002220000022300000224000002250000022600000227),
    .INIT_7D(256'h00002028000002290000022A0000022B0000022C0000022D0000022E0000022F),
    .INIT_7E(256'h0000203000000231000002320000023300000234000002350000023600000237),
    .INIT_7F(256'h00002038000002390000023A0000023B0000023C0000023D0000023E0000023F)

    ) iram_lower (
    .DOA(iram_doa[32:63]),
    .DOB(iram_dob[32:63]),
    .DOPA( ),
    .DOPB( ),
    .ADDRA({1'b0, g_iram_addra, 5'b0}),
    .ADDRB({1'b0, h_iram_addrb, 5'b0}),
    .CLKA(lnk_clk),
    .CLKB(lnk_clk),
    .DIA(32'b0),
    .DIB(32'b0),
    .DIPA(4'b0),
    .DIPB(4'b0),
    .ENA(1'b1),
    .ENB(1'b1),
    .REGCEA(1'b0),
    .REGCEB(1'b0),
    .SSRA(~lnk_reset_n),
    .SSRB(~lnk_reset_n),
    .WEA(4'b0),
    .WEB(4'b0),
    .CASCADEOUTLATA(),
    .CASCADEOUTLATB(),
    .CASCADEOUTREGA(),
    .CASCADEOUTREGB(),
    .CASCADEINLATA(),
    .CASCADEINLATB(),
    .CASCADEINREGA(),
    .CASCADEINREGB()
    );

endmodule
